module ascii_values(Sin,Sout);
input [7:0]Sin;
output [7:0]Sout;
assign Sout=(Sin==8'h45)?8'h30:			//0	100 0000	
		(Sin==8'h16)?8'h31:		//1	111 1001
		(Sin==8'h1E)?8'h32:		//2	010 0100
		(Sin==8'h26)?8'h33:		//3	011 0000
		(Sin==8'h25)?8'h34:		//4	000 1001
		(Sin==8'h2E)?8'h35:		//5	001 0010
		(Sin==8'h36)?8'h36:		//6	000 0010
		(Sin==8'h3D)?8'h37:		//7	111 1000	
		(Sin==8'h3E)?8'h38:		//8	000 0000
		(Sin==8'h46)?8'h39:		//9	001 0000
		(Sin==8'h1C)?8'h41:		//A	000 1000
		(Sin==8'h32)?8'h42:		//b	000 0011
		(Sin==8'h21)?8'h43:		//C	100 0110
		(Sin==8'h23)?8'h44:		//d	010 0001
		(Sin==8'h24)?8'h45:		//E	000 0110
		(Sin==8'h2B)?8'h46:		//F	000 1110
		(Sin==8'h1D)?8'h57:	   
		(Sin==8'h75)?8'h12:8'h2E;	
endmodule
